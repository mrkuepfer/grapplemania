wall 0 0 20 400 white
wall 0 400 20 400 white
wall 0 800 20 400 white
wall 20 1180 400 20 white
wall 420 1180 400 20 white
wall 820 1180 400 20 white
wall 1220 1180 400 20 white
wall 1620 1180 400 20 white
wall 2000 780 20 400 white
wall 2000 380 20 400 white
wall 2000 0 20 380 white
wall 1620 0 380 20 white
wall 1240 0 380 20 white
wall 480 0 380 20 white
wall 20 0 380 20 white
wall 260 0 380 20 white
start 20 20 80 80 green
end 1920 20 80 80 red
wall 360 20 40 500 white
wall 20 720 500 40 white
wall 520 720 300 40 white
wall 780 420 40 300 white
wall 780 140 40 300 white
wall 1140 40 40 300 white
wall 1140 340 40 300 white
wall 1140 640 40 300 white
wall 840 900 300 40 white
wall 540 900 300 40 white
wall 240 900 300 40 white
wall 1440 720 120 120 white
wall 1700 420 120 120 white
wall 1420 160 120 120 white
wall 860 0 380 20 white
