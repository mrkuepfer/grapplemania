wall 0 0 40 520 white
wall 0 520 40 520 white
wall 40 0 520 40 white
wall 560 0 520 40 white
wall 1080 0 40 520 white
wall 1080 520 40 520 white
wall 1080 1040 40 520 white
wall 0 1040 40 520 white
wall 0 1560 40 520 white
wall 1080 1560 40 520 white
wall 0 2080 40 520 white
wall 1080 2080 40 520 white
wall 0 2600 40 520 white
wall 1080 2600 40 520 white
wall 0 3120 40 520 white
wall 1080 3120 40 520 white
wall 1080 3640 40 520 white
wall 0 3640 40 520 white
wall 0 4160 40 520 white
wall 1080 4160 40 520 white
wall 0 4680 40 520 white
wall 1080 4680 40 520 white
wall 0 5200 520 40 white
wall 520 5200 520 40 white
wall 1040 5200 80 40 white
start 540 5160 80 40 green
wall 240 4960 660 40 white
wall 540 4640 40 340 white
wall 540 4320 40 340 white
death 500 4320 40 340 darkmagenta
death 500 4660 40 340 darkmagenta
death 580 4320 40 340 darkmagenta
death 580 4660 40 340 darkmagenta
wall 580 4960 40 40 white
wall 500 4960 40 40 white
death 40 4460 40 400 darkmagenta
death 40 4300 40 160 darkmagenta
death 1040 4320 40 160 darkmagenta
death 1040 4480 40 160 darkmagenta
death 1040 4640 40 160 darkmagenta
death 1040 4800 40 60 darkmagenta
death 160 4120 280 40 darkmagenta
death 700 4120 280 40 darkmagenta
booster 260 4320 40 140 orange
booster 260 4460 40 140 orange
booster 820 4320 40 140 orange
booster 820 4460 40 140 orange
checkpoint 40 3880 1040 40 blue
wall 320 4000 480 40 white
wall 260 3280 40 480 white
wall 540 3280 40 480 white
wall 800 3280 40 480 white
checkpoint 940 3480 40 40 blue
checkpoint 660 3480 40 40 blue
checkpoint 400 3480 40 40 blue
checkpoint 120 3480 40 40 blue
wall 40 3060 800 40 white
wall 280 2740 800 40 white
wall 40 2480 800 40 white
wall 280 2220 800 40 white
booster 140 3020 700 40 orange
booster 280 2700 700 40 orange
booster 140 2440 700 40 orange
booster 280 2180 700 40 orange
death 980 2180 100 40 darkmagenta
death 40 2440 100 40 darkmagenta
death 980 2700 100 40 darkmagenta
death 40 3020 100 40 darkmagenta
checkpoint 40 40 1040 40 blue
wall 20 2020 960 40 white
wall 220 1740 100 100 white
wall 620 1600 100 100 white
wall 380 1420 100 100 white
wall 860 1300 100 100 white
wall 120 1220 100 100 white
wall 580 1120 100 100 white
wall 300 980 100 100 white
wall 820 900 100 100 white
wall 520 720 100 100 white
wall 120 720 100 100 white
wall 800 500 100 100 white
wall 260 280 100 100 white
death 460 480 100 100 darkmagenta
death 380 1180 100 100 darkmagenta
death 980 1080 100 100 darkmagenta
death 40 1560 100 100 darkmagenta
death 980 1480 100 100 darkmagenta
end 540 4996 80 40 red
