wall 0 0 20 400 white
wall 0 400 20 400 white
wall 0 800 20 400 white
wall 20 1180 400 20 white
wall 420 1180 400 20 white
wall 820 1180 400 20 white
wall 1220 1180 400 20 white
wall 1620 1180 400 20 white
wall 2000 780 20 400 white
wall 2000 380 20 400 white
wall 2000 0 20 380 white
wall 1620 0 380 20 white
wall 1240 0 380 20 white
wall 860 0 380 20 white
wall 480 0 380 20 white
wall 20 0 380 20 white
wall 260 0 380 20 white
end 1920 20 80 80 red
wall 20 220 280 40 white
start 20 20 100 200 green
wall 520 20 40 200 white
wall 520 220 40 200 white
wall 360 420 200 40 white
wall 20 620 200 40 white
wall 220 620 200 40 white
wall 420 620 140 40 white
booster 160 520 140 40 orange
booster 300 520 140 40 orange
booster 440 520 120 40 orange
wall 560 620 120 40 white
wall 680 620 120 40 white
wall 760 500 40 120 white
wall 760 380 40 120 white
wall 760 280 40 120 white
wall 760 180 40 120 white
wall 160 420 200 40 white
checkpoint 540 460 20 160 blue
death 740 180 20 160 darkmagenta
death 740 160 80 20 darkmagenta
death 800 180 20 140 darkmagenta
wall 980 20 40 260 white
wall 980 280 40 260 white
wall 980 540 40 260 white
wall 760 800 260 40 white
checkpoint 800 640 180 20 blue
wall 580 800 180 40 white
wall 400 800 180 40 white
wall 220 800 180 40 white
death 660 760 40 40 darkmagenta
death 440 660 40 40 darkmagenta
death 180 800 40 40 darkmagenta
death 20 800 40 40 darkmagenta
wall 220 840 40 160 white
checkpoint 20 980 200 20 blue
wall 440 1100 80 80 white
wall 360 940 80 80 white
wall 560 840 80 80 white
wall 940 840 80 80 white
death 1580 1140 420 40 darkmagenta
death 1960 720 40 420 darkmagenta
death 1960 320 40 420 darkmagenta
death 1020 420 40 420 darkmagenta
death 1020 20 40 400 darkmagenta
death 1060 20 400 40 darkmagenta
death 1460 20 400 40 darkmagenta
death 1960 160 40 160 darkmagenta
wall 734 925 80 80 white
wall 854 1065 80 80 white
wall 1294 725 40 40 white
wall 1734 585 40 40 white
wall 1374 365 40 40 white
wall 1214 165 40 40 white
wall 1654 145 40 40 white
death 800 320 20 20 darkmagenta
